module instruction_memory(rst, addr, ins);
	input rst;
	input [31:0] addr;
	output [31:0] ins;
	reg [31:0] memory[31:0];
		
	always@ (negedge rst) begin
		if (!rst) begin
			//		ADDI	R7, R0, 6
			//		ADDI	R1, R0, 0
			//		ADDI	R2, R0, 1
			//		ADDI	R3, R0, 1
			//		ADDI	R4, R0, 2
			//		J		TES
			//FIB:	ADDI	R4, R4, 1
			//		ADDI	R1, R2, 0
			//		ADDI	R2, R3, 0
			//		ADD	R3, R2, R1
			//		J		OUT
			//TES:	BEQ	R7, R4, OUT
			//		J		FIB
			//OUT:	SW	R3, 0(R0)

			 memory[0] <= 32'b001000_00000_00111_00000_00000_000110;
			 memory[1] <= 32'b001000_00000_00001_00000_00000_000000;
			 memory[2] <= 32'b001000_00000_00010_00000_00000_000001;
			 memory[3] <= 32'b001000_00000_00011_00000_00000_000001;
			 memory[4] <= 32'b001000_00000_00100_00000_00000_000010;
			 memory[5] <= 32'b000010_00000_00000_00000_00001_010000;
			 
			memory[10] <= 32'b001000_00100_00100_00000_00000_000001;
			memory[11] <= 32'b001000_00010_00001_00000_00000_000000;
			memory[12] <= 32'b001000_00011_00010_00000_00000_000000;
			memory[13] <= 32'b000000_00010_00001_00011_00000_100000;
			memory[14] <= 32'b000010_00000_00000_00000_00001_100100;
			
			memory[20] <= 32'b000100_00111_00100_00000_00000_000100;
			memory[21] <= 32'b000010_00000_00000_00000_00000_101000;
			
			memory[25] <= 32'b101011_00000_00011_00000_00000_000000;
			
			memory[31] <= 32'b000000_00000_00000_00000_00000_101001;
			end
	end
	
	assign ins = memory[addr>>2];

endmodule
